library ieee;
use ieee.std_logic_1164.all;

entity andGate is 
	port(
	a , b :in std_logic;
	c : out std_logic
	);
end entity ;

architecture arch of  andGate is 
begin 
	c <= a and b;
	end architecture ;